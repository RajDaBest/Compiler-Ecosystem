#define alloc 0
#define free 1
#define print_f64 2
#define print_s64 3
#define print_u64 4